`timescale 1ns / 1ps
module design_top(

    );
endmodule
