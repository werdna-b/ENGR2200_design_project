`timescale 1ns / 1ps

module counter(
   input enable, clk
   );


endmodule
