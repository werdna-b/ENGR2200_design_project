`timescale 1ns / 1ps


module Lets_go(
    input clk,          // 100 MHz System Clock (Pin W5)
    input mix_state,
    input btnC
    );
    
    always @(posedge clk) begin
    
    
    
    end
    
    
    





endmodule
